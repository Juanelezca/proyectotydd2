library verilog;
use verilog.vl_types.all;
entity control_tiempo_vlg_vec_tst is
end control_tiempo_vlg_vec_tst;
